module conv1_calc_1(
    input valid_out_buf,
    input pixel_0, pixel_1, pixel_2,
        pixel_3, pixel_4, pixel_5,
        pixel_6, pixel_7, pixel_8,
    output reg conv1_out_1, conv1_out_2, conv1_out_3, conv1_out_4,
        conv1_out_5, conv1_out_6, conv1_out_7, conv1_out_8,
    output reg valid_out_conv1
);


endmodule
module conv_layer_2 (
    input wire clk,
    input wire rst_n,
    input wire data_in,         // 1-bit input data
    output reg conv2_out_1,      // 16 channels output signals for convolution layer 2
    output reg conv2_out_2,      // each clk one bit output
    output reg conv2_out_3,
    output reg conv2_out_4,
    output reg conv2_out_5,
    output reg conv2_out_6,
    output reg conv2_out_7,
    output reg conv2_out_8,
    output reg conv2_out_9,
    output reg conv2_out_10,
    output reg conv2_out_11,
    output reg conv2_out_12,
    output reg conv2_out_13,
    output reg conv2_out_14,
    output reg conv2_out_15,
    output reg conv2_out_16,
    output reg valid_out_conv2  // signal to indicate valid output
);


endmodule